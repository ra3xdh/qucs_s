* EF183 Variable-mu Pentode Spice Model
* Author: Zabb Csaba
* Date:   26/10/2021
* The following parameters are not modelled:
*   (1) Filament and filament warmup time
*   (2) Limiting values
.SUBCKT EF183 A S G K 
+ PARAMS: MU=45.58 KG1=126.5 KP=141.9 KVB=12 VCT=6.25E-4 EX=1.008 KG2=258 KNEE=7.92 KVC=2.82
+ KLAM=2E-7 KLAMG=9.9E-5 KNEE2=7.963 KNEX=2.756  
E1  1 0  VALUE={V(S,K)/KP*LOG(1+EXP((1/MU+(VCT+V(G,K)*V(3))/SQRT(KVB+V(S,K)*V(S,K)))*KP))}
E2  2 0  VALUE={(PWR(V(1),EX)+PWRS(V(1),EX))}
G1  A K  VALUE={IF(V(A,K)>0,V(2)/KG1*ATAN((V(A,K)+KNEX)/KNEE)*TANH(V(A,K)/KNEE2)*(1+KLAMG*V(A,K)),0)}
E4  4 K  VALUE={IF(V(A,K)>0,V(A,K),0)}
G2  S K  VALUE={V(2)/KG2*(KVC-ATAN((V(4,K)+KNEX)/KNEE)*TANH(V(4,K)/KNEE2))/(1+KLAMG*V(4,K))}
G3  G K  VALUE={3.16E-2*(PWR(V(G,K),1.5)+PWRS(V(G,K),1.5))/2} ; G1 diode
E3  3 0  VALUE={IF(V(G,K)<0,(1-EXP(14/V(G,K)))^1.3,1)}
B1  G K  I=URAMP(V(G,K)+1.015)^1.5*5.1E-4*V(6)
B2  G K  I=URAMP(V(G,K)+1.015)^1.5*2E-4  
E5  5 0  VALUE={IF(V(S,K)>0,1/(1+ABS(V(S,K))/20)^2,1)} ;G1 Splash current change
E6  6 0  VALUE={IF(V(A,K)>=15,V(5),1)}
C1  G K  9p
C2  A K  3p
C3  A G  0.005p
.ENDS EF183
*$