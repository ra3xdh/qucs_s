*  MOC3063 Zero-Cross Optoisolators Triac Driver Output Spice Model
*  Date  : 08/09/2024
*  Author: Zabb Csaba
*  IRED  emitting  diodes  optically  coupled  to  monolithic  silicon  detectors
*  performing the functions of Zero Voltage Crossing bilateral triac drivers.
*  VINH=Inhibit Voltage (MT1–MT2 Voltage above which device will not trigger.)
*
.SUBCKT MOC3063  1   2   6    4    
*                A   K  MT2  MT1 
DL  1   3   IRLED
V1  3   2   0
H1  17  0   V1  1
E1  DEL 0   TABLE {V(17)}
+ (5m,  50)
+ (10m, 30)
+ (15m, 19)
+ (20m, 14)
+ (25m, 11)
+ (30m, 10)
+ (35m, 9.0)
+ (40m, 8.0)
+ (45m, 7.0)
+ (50m, 6.5)
+ (55m, 6.1)
E2  11  0   VALUE {IF(V(17)>5m,1,0)}
X1  11  10  DEL 0 VCRES
C1  10  0   1n
E3  12  4   VALUE {IF(V(10)>0.63,1,0)}
S1  6   13  11  0 SW1
R1  13  8   3MEG
C2  8   4   10p
D1  8   7   DX
D2  4   7   DX 
E4  9   4   VALUE {IF(ABS(V(8,4))<12,1,0)}
B1  G   4   I=V(12,4)*V(9,4)*10m
C3  2   4   800f
R2  2   4   10G
X2  6   4   G   TRIAC Ih=0.25m
.MODEL  DX D(BV=50 IBV=10u)
.MODEL  SW1 VSWITCH (ROFF=1G RON=1 VOFF=0 VON=1)
.MODEL  IRLED D (IS=8E-17 N=1.5 RS=2 IKF=7.5E-2 IBV=1.5E-08 NBV=7E1  BV=1.6E1 CJO=4E-11 TT=1E-08 EG=1.46)
.ENDS MOC3063

*  Author: Zabb Csaba
*  IRED emitting diode optically coupled to a non-zero-crossing silicon bilateral AC switch (triac).
*
.SUBCKT MOC3052  1   2   6    4   
*                A   K  MT2  MT1 
DL  1   5   IRLED
V1  5   2   0
H1  7   0   V1  1
E1  DEL 0   TABLE {V(7)}
+ (10m, 30)
+ (15m, 19)
+ (20m, 14)
+ (25m, 11)
+ (30m, 10)
+ (35m, 9.0)
+ (40m, 8.0)
+ (45m, 7.0)
+ (50m, 6.5)
+ (55m, 6.1)
E2  11  0   VALUE {IF(V(7)>10m,1,0)}
X1  11  9   DEL 0 VCRES
C1  9   0   1n
E3  8   4   VALUE {IF(V(9)>0.63,1,0)}
G1  G   4   8   4   10m
C2  2   4   800f
R1  2   4   10G
X2  6   4   G   TRIAC Ih=0.28m
.MODEL  IRLED D (IS=8E-17 N=1.5 RS=2 IKF=7.5E-2 IBV=1.5E-08 NBV=7E1 BV=1.6E1 CJO=4E-11 TT=1E-08 EG=1.46)
.ENDS MOC3052

*
.SUBCKT VCRES	1 2	4 5
+PARAMS: R1=1k
ERES	1	3	VALUE={IF(V(4,5)>0,I(VSENSE)*{R1}*V(4,5),-I(VSENSE)*{R1}*V(4,5))}
VSENSE	3	2	0
.ENDS VCRES
*
.SUBCKT TRIAC MT2 MT1 G params:
+ Vdrm=600   
+ Igt=5m
+ Ih=0.28m       
+ Rt=3.3
+ Standard=1
S1  MT2 2   3   0 SW1
D1  2   4   DAK 
R1  2   4   1k
V1  4   MT1 0
S2  MT2 5   6   0 SW1
D2  7   5   DAK 
R2  5   7   1k 
V2  MT1 7   0 
R3  G   MT1 1G  
D3  8   G   DGK 
D4  G   8   DGK 
V3  8   MT1 0 
R4  G   8   1k  
R5  9   3   2.2  
C1  0   3   5u 
E1  9   0   VALUE {IF(((V(10)>0.5)|(V(13)>0.5)|(V(12)>0.5)),400,0)}
R6  14  6   2.2   
C2  0   6   5u  
E2  14  0   VALUE {IF(((V(10)>0.5)|(V(11)>0.5)|(V(12)>0.5)),400,0)}
E3  15  0   VALUE {IF((ABS(I(V3)))>(Igt-1u),1,0)}
E4  16  0   VALUE {V(17)*V(15)}
E5  17  0   VALUE {IF(((I(V3)>(Igt-1u))&((V(MT2)-V(MT1))<0)&(Standard==0)),0,1)}
X1  16  10  BUFDELAY
E6  18  0   VALUE {IF(((I(V1))>(Ih/2)),1,0)}
E7  19  0   VALUE {IF(((I(V1))>(Ih/3)),1,0)} 
E8  20  0   VALUE {IF((V(18)*V(19)+V(19)*(1-V(18))*(V(21)))>0.5,1,0)}
C3  21  0   1n  
R7  20  21  1k  
R8  21  0   100MEG  
X2  21  13  BUFDELAY
E9  22  0   VALUE {IF(((I(V2))>(Ih/2)),1,0)}
E10 23  0   VALUE {IF(((I(V2))>(Ih/3)),1,0)} 
E11 24  0   VALUE {IF((V(22)*V(23)+V(23)*(1-V(22))*(V(25)))>0.5,1,0)}
C4  25  0   1n  
R9  24  25  1k  
R10 25  0   100MEG 
X3  25  11  BUFDELAY
E12 26  0   VALUE {IF((ABS(V(MT2)-V(MT1))>(Vdrm*1.3)),1,0)}
E13 27  0   VALUE {IF((I(V1)>(Vdrm*1.3)/5MEG)|(I(V2)>(Vdrm*1.3)/5MEG),1,0)}
E14 28  0   VALUE {IF((V(26)+(1-V(26))*V(27)*V(29) )>0.5,1,0)}
C5  29  0   1n  
R11 28  29  100  
R12 29  0   100MEG 
X4  29  12  BUFDELAY
.MODEL  SW1 VSWITCH (ROFF=1G RON={Rt} VOFF=0 VON=1)
.MODEL  DAK D(IS=3E-12 N=1.66 CJO=5p) 
.MODEL  DGK D(IS=1E-16 CJO=50p Rs=5) 
.ENDS TRIAC
*
.SUBCKT BUFDELAY A Y PARAMS:DELAY=1u 
E1 Y1 0  VALUE {IF(V(A)>0.5,1,0)}
R1 Y1 Y2 1
C1 Y2 0  {DELAY*1.44}
E2 Y3 0  VALUE {IF(V(Y2)>0.5,1,0)}
R2 Y3 Y  1
C2 Y  0  1n
.ENDS BUFDELAY
*$