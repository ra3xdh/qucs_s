* 6K1J Variable-mu VHF Pentode Spice Model
* Author: Zabb Csaba
* Date:   6/11/2021
* The following parameters are not modelled:
*   (1) Filament and filament warmup time
*   (2) Limiting values
* This model is valid for the following tubes (within max. ratings):
* RCA 956, VT-238, E2F
.SUBCKT 6K1J A S G K 
+ PARAMS: MU=19.2 KG1=95744 KP=12.95 KVB=5.76 VCT=0.0575 EX=2.828 KG2=120960 KNEE=14.4 KVC=2.339
+ KLAM=2.5E-8 KLAMG=7.8E-5 KNEE2=13.39 KNEX=11.1  
E1 1 0  VALUE={V(S,K)/KP*LOG(1+EXP((1/MU+(VCT+V(G,K)*V(3))/SQRT(KVB+V(S,K)*V(S,K)))*KP))}
E3 3 0  VALUE={ATAN(V(G,K)/19+1)/2.7+0.5}
E2 2 0  VALUE={(PWR(V(1),EX)+PWRS(V(1),EX))}
G1 A K  VALUE={IF(V(A,K)>0,0.831*V(2)/KG1*ATAN((V(A,K)+KNEX)/KNEE)*TANH(V(A,K)/KNEE2)*(1+KLAMG*V(A,K)),0)}
E4 4 K  VALUE={IF(V(A,K)>0,V(A,K),0)}
G2 S K  VALUE={0.822*V(2)/KG2*(KVC-ATAN((V(4,K)+KNEX)/KNEE)*TANH(V(4,K)/KNEE2))/(1+KLAMG*V(4,K))}
B1 G K  I=URAMP(V(G,K)+1.15)^1.5*2.6E-4*V(5)
E5 5 0  VALUE={IF(V(S,K)>0,1/(1+ABS(V(S,K))/20)^1.3,1)} ;G1 Splash current change
R1 5 0  1G
C1 G K  3.4p
C2 A K  3p
C3 G A  0.007p
.ENDS
*$